module sbox(byte_in, byte_out, clk);

  input [7:0] byte_in;
  output [7:0] byte_out;
  input clk;

  reg [7:0] byte_out;
  reg [7:0] rom [0:255];

  initial begin
    rom[  0] <= 8'h63;
    rom[  1] <= 8'h7C;
    rom[  2] <= 8'h77;
    rom[  3] <= 8'h7B;
    rom[  4] <= 8'hF2;
    rom[  5] <= 8'h6B;
    rom[  6] <= 8'h6F;
    rom[  7] <= 8'hC5;
    rom[  8] <= 8'h30;
    rom[  9] <= 8'h01;
    rom[ 10] <= 8'h67;
    rom[ 11] <= 8'h2B;
    rom[ 12] <= 8'hFE;
    rom[ 13] <= 8'hD7;
    rom[ 14] <= 8'hAB;
    rom[ 15] <= 8'h76;
    rom[ 16] <= 8'hCA;
    rom[ 17] <= 8'h82;
    rom[ 18] <= 8'hC9;
    rom[ 19] <= 8'h7D;
    rom[ 20] <= 8'hFA;
    rom[ 21] <= 8'h59;
    rom[ 22] <= 8'h47;
    rom[ 23] <= 8'hF0;
    rom[ 24] <= 8'hAD;
    rom[ 25] <= 8'hD4;
    rom[ 26] <= 8'hA2;
    rom[ 27] <= 8'hAF;
    rom[ 28] <= 8'h9C;
    rom[ 29] <= 8'hA4;
    rom[ 30] <= 8'h72;
    rom[ 31] <= 8'hC0;
    rom[ 32] <= 8'hB7;
    rom[ 33] <= 8'hFD;
    rom[ 34] <= 8'h93;
    rom[ 35] <= 8'h26;
    rom[ 36] <= 8'h36;
    rom[ 37] <= 8'h3F;
    rom[ 38] <= 8'hF7;
    rom[ 39] <= 8'hCC;
    rom[ 40] <= 8'h34;
    rom[ 41] <= 8'hA5;
    rom[ 42] <= 8'hE5;
    rom[ 43] <= 8'hF1;
    rom[ 44] <= 8'h71;
    rom[ 45] <= 8'hD8;
    rom[ 46] <= 8'h31;
    rom[ 47] <= 8'h15;
    rom[ 48] <= 8'h04;
    rom[ 49] <= 8'hC7;
    rom[ 50] <= 8'h23;
    rom[ 51] <= 8'hC3;
    rom[ 52] <= 8'h18;
    rom[ 53] <= 8'h96;
    rom[ 54] <= 8'h05;
    rom[ 55] <= 8'h9A;
    rom[ 56] <= 8'h07;
    rom[ 57] <= 8'h12;
    rom[ 58] <= 8'h80;
    rom[ 59] <= 8'hE2;
    rom[ 60] <= 8'hEB;
    rom[ 61] <= 8'h27;
    rom[ 62] <= 8'hB2;
    rom[ 63] <= 8'h75;
    rom[ 64] <= 8'h09;
    rom[ 65] <= 8'h83;
    rom[ 66] <= 8'h2C;
    rom[ 67] <= 8'h1A;
    rom[ 68] <= 8'h1B;
    rom[ 69] <= 8'h6E;
    rom[ 70] <= 8'h5A;
    rom[ 71] <= 8'hA0;
    rom[ 72] <= 8'h52;
    rom[ 73] <= 8'h3B;
    rom[ 74] <= 8'hD6;
    rom[ 75] <= 8'hB3;
    rom[ 76] <= 8'h29;
    rom[ 77] <= 8'hE3;
    rom[ 78] <= 8'h2F;
    rom[ 79] <= 8'h84;
    rom[ 80] <= 8'h53;
    rom[ 81] <= 8'hD1;
    rom[ 82] <= 8'h00;
    rom[ 83] <= 8'hED;
    rom[ 84] <= 8'h20;
    rom[ 85] <= 8'hFC;
    rom[ 86] <= 8'hB1;
    rom[ 87] <= 8'h5B;
    rom[ 88] <= 8'h6A;
    rom[ 89] <= 8'hCB;
    rom[ 90] <= 8'hBE;
    rom[ 91] <= 8'h39;
    rom[ 92] <= 8'h4A;
    rom[ 93] <= 8'h4C;
    rom[ 94] <= 8'h58;
    rom[ 95] <= 8'hCF;
    rom[ 96] <= 8'hD0;
    rom[ 97] <= 8'hEF;
    rom[ 98] <= 8'hAA;
    rom[ 99] <= 8'hFB;
    rom[100] <= 8'h43;
    rom[101] <= 8'h4D;
    rom[102] <= 8'h33;
    rom[103] <= 8'h85;
    rom[104] <= 8'h45;
    rom[105] <= 8'hF9;
    rom[106] <= 8'h02;
    rom[107] <= 8'h7F;
    rom[108] <= 8'h50;
    rom[109] <= 8'h3C;
    rom[110] <= 8'h9F;
    rom[111] <= 8'hA8;
    rom[112] <= 8'h51;
    rom[113] <= 8'hA3;
    rom[114] <= 8'h40;
    rom[115] <= 8'h8F;
    rom[116] <= 8'h92;
    rom[117] <= 8'h9D;
    rom[118] <= 8'h38;
    rom[119] <= 8'hF5;
    rom[120] <= 8'hBC;
    rom[121] <= 8'hB6;
    rom[122] <= 8'hDA;
    rom[123] <= 8'h21;
    rom[124] <= 8'h10;
    rom[125] <= 8'hFF;
    rom[126] <= 8'hF3;
    rom[127] <= 8'hD2;
    rom[128] <= 8'hCD;
    rom[129] <= 8'h0C;
    rom[130] <= 8'h13;
    rom[131] <= 8'hEC;
    rom[132] <= 8'h5F;
    rom[133] <= 8'h97;
    rom[134] <= 8'h44;
    rom[135] <= 8'h17;
    rom[136] <= 8'hC4;
    rom[137] <= 8'hA7;
    rom[138] <= 8'h7E;
    rom[139] <= 8'h3D;
    rom[140] <= 8'h64;
    rom[141] <= 8'h5D;
    rom[142] <= 8'h19;
    rom[143] <= 8'h73;
    rom[144] <= 8'h60;
    rom[145] <= 8'h81;
    rom[146] <= 8'h4F;
    rom[147] <= 8'hDC;
    rom[148] <= 8'h22;
    rom[149] <= 8'h2A;
    rom[150] <= 8'h90;
    rom[151] <= 8'h88;
    rom[152] <= 8'h46;
    rom[153] <= 8'hEE;
    rom[154] <= 8'hB8;
    rom[155] <= 8'h14;
    rom[156] <= 8'hDE;
    rom[157] <= 8'h5E;
    rom[158] <= 8'h0B;
    rom[159] <= 8'hDB;
    rom[160] <= 8'hE0;
    rom[161] <= 8'h32;
    rom[162] <= 8'h3A;
    rom[163] <= 8'h0A;
    rom[164] <= 8'h49;
    rom[165] <= 8'h06;
    rom[166] <= 8'h24;
    rom[167] <= 8'h5C;
    rom[168] <= 8'hC2;
    rom[169] <= 8'hD3;
    rom[170] <= 8'hAC;
    rom[171] <= 8'h62;
    rom[172] <= 8'h91;
    rom[173] <= 8'h95;
    rom[174] <= 8'hE4;
    rom[175] <= 8'h79;
    rom[176] <= 8'hE7;
    rom[177] <= 8'hC8;
    rom[178] <= 8'h37;
    rom[179] <= 8'h6D;
    rom[180] <= 8'h8D;
    rom[181] <= 8'hD5;
    rom[182] <= 8'h4E;
    rom[183] <= 8'hA9;
    rom[184] <= 8'h6C;
    rom[185] <= 8'h56;
    rom[186] <= 8'hF4;
    rom[187] <= 8'hEA;
    rom[188] <= 8'h65;
    rom[189] <= 8'h7A;
    rom[190] <= 8'hAE;
    rom[191] <= 8'h08;
    rom[192] <= 8'hBA;
    rom[193] <= 8'h78;
    rom[194] <= 8'h25;
    rom[195] <= 8'h2E;
    rom[196] <= 8'h1C;
    rom[197] <= 8'hA6;
    rom[198] <= 8'hB4;
    rom[199] <= 8'hC6;
    rom[200] <= 8'hE8;
    rom[201] <= 8'hDD;
    rom[202] <= 8'h74;
    rom[203] <= 8'h1F;
    rom[204] <= 8'h4B;
    rom[205] <= 8'hBD;
    rom[206] <= 8'h8B;
    rom[207] <= 8'h8A;
    rom[208] <= 8'h70;
    rom[209] <= 8'h3E;
    rom[210] <= 8'hB5;
    rom[211] <= 8'h66;
    rom[212] <= 8'h48;
    rom[213] <= 8'h03;
    rom[214] <= 8'hF6;
    rom[215] <= 8'h0E;
    rom[216] <= 8'h61;
    rom[217] <= 8'h35;
    rom[218] <= 8'h57;
    rom[219] <= 8'hB9;
    rom[220] <= 8'h86;
    rom[221] <= 8'hC1;
    rom[222] <= 8'h1D;
    rom[223] <= 8'h9E;
    rom[224] <= 8'hE1;
    rom[225] <= 8'hF8;
    rom[226] <= 8'h98;
    rom[227] <= 8'h11;
    rom[228] <= 8'h69;
    rom[229] <= 8'hD9;
    rom[230] <= 8'h8E;
    rom[231] <= 8'h94;
    rom[232] <= 8'h9B;
    rom[233] <= 8'h1E;
    rom[234] <= 8'h87;
    rom[235] <= 8'hE9;
    rom[236] <= 8'hCE;
    rom[237] <= 8'h55;
    rom[238] <= 8'h28;
    rom[239] <= 8'hDF;
    rom[240] <= 8'h8C;
    rom[241] <= 8'hA1;
    rom[242] <= 8'h89;
    rom[243] <= 8'h0D;
    rom[244] <= 8'hBF;
    rom[245] <= 8'hE6;
    rom[246] <= 8'h42;
    rom[247] <= 8'h68;
    rom[248] <= 8'h41;
    rom[249] <= 8'h99;
    rom[250] <= 8'h2D;
    rom[251] <= 8'h0F;
    rom[252] <= 8'hB0;
    rom[253] <= 8'h54;
    rom[254] <= 8'hBB;
    rom[255] <= 8'h16;
  end

  always @(posedge clk) begin
      byte_out <= rom[byte_in];
  end
endmodule


